`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:51:27 02/21/2018 
// Design Name: 
// Module Name:    instruction 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module instruction(input [31:0] readAdd,
						 output reg [31:0] out
    );
	
	always @(*)
		case(readAdd)
			32'b0: out = 32'b000000_00000_00001_00010_00000_100000; // 1+2=3  3 to reg 2
			32'b1: out = 32'b000000_00000_00001_00010_00000_100010; // 1-2=-1 to reg2
			32'b10: out = 32'b000000_00000_00001_00010_00000_100100; //and
			32'b11: out = 32'b000000_00000_00001_00010_00000_100101; //or
			32'b100: out = 32'b000000_00000_00001_00010_00000_100100; //and			
			32'b101: out = 32'b000010_00000000000000000000001000;//jump to add pc+2
			
			32'b110: out = 32'b101011_00100_00011_0000000000000101;//store 5 to mem 3
			32'b111: out = 32'b100011_00100_00011_00000000000000100;//load 4 in reg 3
			
			32'b1000: out = 32'b000000_00000_00001_00010_00000_100000; // 1+2=3  3 to reg 2
    		32'b1001: out = 32'b000000_00000_00001_00010_00000_100010; // 1-2=-1 to reg2
		   32'b1010: out = 32'b000000_00000_00001_00010_00000_100100; //and
			32'b1011: out = 32'b000000_00000_00001_00010_00000_100101; //or
			
			default: out = 32'b00000000000000000000000000000000;
		endcase
endmodule
